/*
 * Copyright (C) 2010, Jason S. McMullan. All rights reserved.
 * Author: Jason S. McMullan <jason.mcmullan@gmail.com>
 *
 * This program is free software; you can redistribute it and/or
 * modify it under the terms of the GNU General Public License
 * as published by the Free Software Foundation; either version 2
 * of the License, or (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with this program; if not, write to the Free Software
 * Foundation, Inc., 51 Franklin Street, Fifth Floor,
 * Boston, MA 02110-1301, USA.
 *
 */

module RAM_41464 (
	input	_OE,
	inout	DQ1,
	inout	DQ2,
	input	_W,
	input	_RAS,
	input	A6,
	input	A5,
	input	A4,
	input	VCC,
	input	A7,
	input	A3,
	input	A2,
	input	A1,
	input	A0,
	inout	DQ3,
	input	_CAS,
	inout	DQ4,
	input	GND
);

// TODO: Implement this!

endmodule
